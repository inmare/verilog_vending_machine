`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/12/03 20:17:23
// Design Name: 
// Module Name: item_based_piezo
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module item_based_piezo(
    input clk, rst,
    input [3:0] note_state,
    input [2:0] note_played,
    output reg piezo
    );

    // piezo�� ���̸� ���ļ�
    reg [11:0] piezo_limit;
    parameter xx = 12'd0;
    parameter do = 12'd3830;
    parameter re = 12'd3400;
    parameter mi = 12'd3038;
    parameter fa = 12'd2864;
    parameter so = 12'd2550;
    parameter la = 12'd2272;
    parameter ti = 12'd2028;
    parameter high_do = 12'd1912;

    parameter note_100w = 1;
    parameter note_500w = 2;
    parameter note_1000w = 3;
    parameter note_prod1 = 4;
    parameter note_prod2 = 5;
    parameter note_prod3 = 6;
    parameter note_prod4 = 7;

    parameter [12*4-1:0] note_100w_lut = { do, mi, so, so };
    parameter [12*4-1:0] note_500w_lut = { re, fa, la, la };
    parameter [12*4-1:0] note_1000w_lut = { mi, so, ti, ti };
    parameter [12*4-1:0] note_prod1_lut = { do, xx, do, xx };
    parameter [12*4-1:0] note_prod2_lut = { re, xx, re, xx };
    parameter [12*4-1:0] note_prod3_lut = { mi, xx, mi, xx };
    parameter [12*4-1:0] note_prod4_lut = { fa, xx, fa, xx };

    // ��Ʈ�� �����ϴ� always��
    always @(negedge rst, posedge clk) begin
        if (!rst) begin
            piezo_limit = xx;
        end
        else begin
            // ��Ʈ ī���͸� 1�� �����ϰ� Ư�� ���� ������ ��Ʈ ���� ���¸� ��Ȱ��ȭ �ϰ� ī���͸� �ʱ�ȭ
            case (note_played)
                1 : begin
                    case (note_state)
                        note_100w : piezo_limit = note_100w_lut[12*4-1:12*3];
                        note_500w : piezo_limit = note_500w_lut[12*4-1:12*3];
                        note_1000w : piezo_limit = note_1000w_lut[12*4-1:12*3];
                        note_prod1 : piezo_limit = note_prod1_lut[12*4-1:12*3];
                        note_prod2 : piezo_limit = note_prod2_lut[12*4-1:12*3];
                        note_prod3 : piezo_limit = note_prod3_lut[12*4-1:12*3];
                        note_prod4 : piezo_limit = note_prod4_lut[12*4-1:12*3];
                        default : piezo_limit = xx;
                    endcase
                end
                2 : begin
                    case (note_state)
                        note_100w : piezo_limit = note_100w_lut[12*3-1:12*2];
                        note_500w : piezo_limit = note_500w_lut[12*3-1:12*2];
                        note_1000w : piezo_limit = note_1000w_lut[12*3-1:12*2];
                        note_prod1 : piezo_limit = note_prod1_lut[12*3-1:12*2];
                        note_prod2 : piezo_limit = note_prod2_lut[12*3-1:12*2];
                        note_prod3 : piezo_limit = note_prod3_lut[12*3-1:12*2];
                        note_prod4 : piezo_limit = note_prod4_lut[12*3-1:12*2];
                        default : piezo_limit = xx;
                    endcase
                end
                3 : begin
                    case (note_state)
                        note_100w : piezo_limit = note_100w_lut[12*2-1:12*1];
                        note_500w : piezo_limit = note_500w_lut[12*2-1:12*1];
                        note_1000w : piezo_limit = note_1000w_lut[12*2-1:12*1];
                        note_prod1 : piezo_limit = note_prod1_lut[12*2-1:12*1];
                        note_prod2 : piezo_limit = note_prod2_lut[12*2-1:12*1];
                        note_prod3 : piezo_limit = note_prod3_lut[12*2-1:12*1];
                        note_prod4 : piezo_limit = note_prod4_lut[12*2-1:12*1];
                        default : piezo_limit = xx;
                    endcase
                end
                4 : begin
                    case (note_state)
                        note_100w : piezo_limit = note_100w_lut[12*1-1:12*0];
                        note_500w : piezo_limit = note_500w_lut[12*1-1:12*0];
                        note_1000w : piezo_limit = note_1000w_lut[12*1-1:12*0];
                        note_prod1 : piezo_limit = note_prod1_lut[12*1-1:12*0];
                        note_prod2 : piezo_limit = note_prod2_lut[12*1-1:12*0];
                        note_prod3 : piezo_limit = note_prod3_lut[12*1-1:12*0];
                        note_prod4 : piezo_limit = note_prod4_lut[12*1-1:12*0];
                        default : piezo_limit = xx;
                    endcase
                end
                default : begin
                    piezo_limit = xx;
                end
            endcase
        end
    end

    // piezo�� ī����
    integer piezo_cnt;
    always @(negedge rst, posedge clk) begin
        if (!rst) begin
            piezo <= 0;
            piezo_cnt <= 0;
        end 
        else if (piezo_cnt >= piezo_limit/2) begin
            piezo <= ~piezo;
            piezo_cnt <= 0;
        end
        else piezo_cnt <= piezo_cnt + 1;
    end
endmodule
