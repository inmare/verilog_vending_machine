`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/12/06 09:43:49
// Design Name: 
// Module Name: prod_based_led
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module prod_based_led(
    input clk, rst,
    input [3:0] prod_count_current,
    output reg [3:0] cled_r, cled_g, cled_b
    );
endmodule
