`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/12/03 15:50:30
// Design Name: 
// Module Name: main_logic
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module main_logic(
    input clk, rst,
    input [11:0] button_sw,
    // ���������� fnd array�� ǥ�õ� ��
    output reg [7:0] display_money_binary,
    // text lcd�� ���� ��ǰ ����
    output reg [2:0] prod1_count, prod2_count, prod3_count,
    // piezo�� ���� ������ ��ǰ
    output reg [2:0] selected_item,
    // line1, line2�� ����� ���ڿ��� �����ϴ� ����
    output reg [8*16-1:0] line1_text, line2_text,
    // Ŀ�� �ּҸ� �����ϴ� ����
    output reg [6:0] ddram_address
    );
    // generate���� ����
    genvar i;
    // ���� �Է��� �ݾ��� �����ֱ� ���� cnt
    // ���� ���� 2000000���� �����ؾ� ��
    integer coin_btn_cnt;
    // parameter coin_btn_cnt_limit = 20;
    parameter coin_btn_cnt_limit = 2000000;

    // �ݾ� ��ȯ�� �ݾ��� �����ֱ� ���� cnt
    // ���� ���� 1000000���� �����ؾ� ��
    integer return_cnt;
    // parameter return_cnt_limit = 10;
    parameter return_cnt_limit = 1000000;

    // Ŀ�� �̵� ��ư
    wire move_up_sw, move_down_sw;
    one_shot_en_sw move_up(
        .clk(clk),
        .enable(button_sw[10]),
        .eout(move_up_sw)
    );
    one_shot_en_sw move_down(
        .clk(clk),
        .enable(button_sw[4]),
        .eout(move_down_sw)
    );  

    wire select_toggle_sw;
    // ���� ��ư
    one_shot_en_sw select_toggle(
        .clk(clk),
        .enable(button_sw[7]),
        .eout(select_toggle_sw)
    );

    // ���� �Է� ����ġ
    wire [2:0] coin_btn_sw;
    generate
        for (i = 0; i < 3; i = i + 1) begin
            one_shot_en_sw coin_btn(
                .clk(clk),
                .enable(button_sw[i]),
                .eout(coin_btn_sw[i])
            );
        end
    endgenerate

    // ���� ����ġ
    wire buy_sw;
    one_shot_en_sw buy(
        .clk(clk),
        .enable(button_sw[9]),
        .eout(buy_sw)
    );

    // ��ȯ ����ġ
    wire return_sw;
    one_shot_en_sw return(
        .clk(clk),
        .enable(button_sw[3]),
        .eout(return_sw)
    );

    // �� ��ǰ id
    parameter prod1_id = 1;
    parameter prod2_id = 2;
    parameter prod3_id = 3;

    // �� ��ǰ ����
    parameter prod1_price = 10;
    parameter prod2_price = 12;
    parameter prod3_price = 15;

    // �� ��ǰ �ʱ� ����
    parameter prod1_init_count = 4;
    parameter prod2_init_count = 1;
    parameter prod3_init_count = 0;

    // ���� Ŀ�� ��ġ
    reg [2:0] cursor_pos;
    // ����, �̼��� ����
    reg selected;

    // ���� �Էµ� ��
    reg [7:0] inserted_money;

    // ��� �����丮 ���� ����� �� 10���� ���� ���� ����
    reg [7*9-1:0] total_money_history;
    reg history_disabled;

    // ���� �Է� ����ġ�� ���������� �˷��ִ� state
    reg coin_btn_state;
    // ��ȯ ����ġ�� ���������� �˷��ִ� state
    reg return_state;

    // ��ǰ���� �����ϴ� ����
    // �ִ� 5����, 3���� ��ǰ���� ����
    parameter [8*7*3-1:0] product = {
        // "1.Coke "
        8'h31, 8'h2e, 8'h43, 8'h6f, 8'h6b, 8'h65, 8'h20,
        // "2.Water"
        8'h32, 8'h2e, 8'h57, 8'h61, 8'h74, 8'h65, 8'h72,
        // "3.Juice"
        8'h33, 8'h2e, 8'h4a, 8'h75, 8'h69, 8'h63, 8'h65
        };

    // ������ ���ڷ� �ٲ㼭 �����ϴ� ����
    // 100�� ������ ������ �����ϱ� ������ 100���� ���� ���� ����
    // ���� 2���ڸ� ������ ��
    parameter [8*2*3-1:0] price_text = {
        8'h31, 8'h30, // "10"
        8'h31, 8'h32, // "12"
        8'h31, 8'h35  // "15"
        };

    // ���� lcd�� ǥ�õ� ��ǰ�� ǥ���ϴ� ����
    reg [2:0] line1_prod, line2_prod;

    // ���� ���Ž� �ݾ� ��ȭ�� always��
    always @(negedge rst, posedge clk) begin
        if (!rst) begin
            // ���� ���� �ʱ�ȭ
            selected_item <= 0;
            cursor_pos <= 0;
            selected <= 0;
            inserted_money <= 0;
            total_money_history <= 0;
            prod1_count <= prod1_init_count;
            prod2_count <= prod2_init_count;
            prod3_count <= prod3_init_count;
            coin_btn_state <= 0;
            return_state <= 0;
            history_disabled <= 0;
            coin_btn_cnt <= 0;
            return_cnt <= 0;
            display_money_binary <= 0;
            line1_text <= 0;
            line2_text <= 0;
            ddram_address <= 7'hd;
            // "1.Coke  1000W  ^"
            line1_text[8*16-1:8*9] <= product[8*7*3-1:8*7*2]; // "1.Coke "
            line1_text[8*9-1:8*8] <= 8'h20; // space
            line1_text[8*8-1:8*6] <= price_text[8*2*3-1:8*2*2]; // "10"
            line1_text[8*6-1:8*0] <= {8'h30, 8'h30, 8'h57, 8'h20, 8'h20, 8'h5e}; // "00W  ^"
            // "2.Water 1200W  v"
            line2_text[8*16-1:8*9] <= product[8*7*2-1:8*7*1]; // "2.Water"
            line2_text[8*9-1:8*8] <= 8'h20; // space
            line2_text[8*8-1:8*6] <= price_text[8*2*2-1:8*2*1]; // "12"
            line2_text[8*6-1:8*0] <= {8'h30, 8'h30, 8'h57, 8'h20, 8'h20, 8'h76}; // "00W  v"
        end
        else begin
            // move up ��ư�� ������ ��� Ŀ�� ��ġ�� �� ĭ ���� �̵�
            if (move_up_sw) begin
                if (cursor_pos > 0) begin
                    cursor_pos = cursor_pos - 1;
                    ddram_address = 7'hd;
                end
            end
            // move down ��ư�� ������ ��� Ŀ�� ��ġ�� �� ĭ �Ʒ��� �̵�
            else if (move_down_sw) begin
                if (cursor_pos < 2) begin
                    cursor_pos = cursor_pos + 1;
                    ddram_address = 7'h4d;
                end
            end
            // ���� ��ư�� ������ ���
            else if (select_toggle_sw) begin
                // ������ ������ id�� cursor ��ġ�� + 1�� �� ������ ������
                if (selected_item != 0 && cursor_pos + 1 == selected_item) begin
                    selected_item = 0;
                    selected = 0;
                end
                else begin
                    case (cursor_pos)
                        0 : begin
                            if (prod1_count != 0) begin
                                selected_item = prod1_id;
                                selected = 1;
                            end 
                            // else begin
                            //     selected_item = 0;
                            //     selected = 0;
                            // end
                        end
                        1 : begin
                            if (prod2_count != 0) begin
                                selected_item = prod2_id;
                                selected = 1;
                            end 
                            // else begin
                            //     selected_item = 0;
                            //     selected = 0;
                            // end
                        end
                        2 : begin
                            if (prod3_count != 0) begin
                                selected_item = prod3_id;
                                selected = 1;
                            end 
                            // else begin
                            //     selected_item = 0;
                            //     selected = 0;
                            // end
                        end
                        default : selected_item = 0;
                    endcase
                end
            end
            // ���� �Է� ����ġ�� ������ ��
            else if (coin_btn_sw != 0) begin
                // ��ư ����ġ�� ���� inserted_money�� �ݾ��� ����
                case (coin_btn_sw)
                    3'b100: inserted_money = 1;
                    3'b010: inserted_money = 5;
                    3'b001: inserted_money = 10;
                    default: inserted_money = 0;
                endcase
                // �� �Է� �ݾ� ���縦 �� ĭ�� �ڷ� �а�, 
                // ���� �ֱ� �Է� �ݾ��� �߰��� ���� �迭 ���� �տ� ����
                total_money_history[7*8-1:0] = total_money_history[7*9-1:7*1];
                total_money_history[7*9-1:7*8] = total_money_history[7*8-1:7*7] + inserted_money;
                // ǥ�õǴ� ���� ���Ե� ������ ����
                display_money_binary = inserted_money;
                // ���� �Է� state Ȱ��ȭ
                coin_btn_state = 1;
            end
            // ���� ����ġ�� ������ ��
            else if (buy_sw) begin
                // ���� ������ ��ǰ�� ����
                case (selected_item)
                    prod1_id: begin
                        // ��ī�ݶ��� ������ 0���� ũ�� �� �ݾ��� ��ī�ݶ��� ���ݺ��� ũ��
                        if (prod1_count > 0 && total_money_history[7*9-1:7*8] > prod1_price) begin
                            // ��ī�ݶ��� ������ �ϳ� ���̰�
                            prod1_count = prod1_count - 1;
                            // ��ī�ݶ��� ���ݸ�ŭ �� �ݾ��� ���δ�
                            total_money_history[7*9-1:7*8] = total_money_history[7*9-1:7*8] - prod1_price;
                            // �� �ݾ� ���縦 ���� �ֱ� ���縦 �����ϰ� ���� �ʱ�ȭ
                            total_money_history[7*8-1:7*0] = 0;
                            // ���� �ʱ�ȭ ���� Ȱ��ȭ
                            history_disabled = 1;
                            // ������ ��ǰ�� ���� ���θ� �ʱ�ȭ
                            selected_item = 0;
                            selected = 0;
                        end
                    end
                    prod2_id: begin
                        if (prod2_count > 0 && total_money_history[7*9-1:7*8] > prod2_price) begin
                            prod2_count = prod2_count - 1;
                            total_money_history[7*9-1:7*8] = total_money_history[7*9-1:7*8] - prod2_price;
                            total_money_history[7*8-1:7*0] = 0;
                            history_disabled = 1;
                            selected_item = 0;
                            selected = 0;
                        end
                    end
                    prod3_id: begin
                        if (prod3_count > 0 && total_money_history[7*9-1:7*8] > prod3_price) begin
                            prod3_count = prod3_count - 1;
                            total_money_history[7*9-1:7*8] = total_money_history[7*9-1:7*8] - prod3_price;
                            total_money_history[7*8-1:7*0] = 0;
                            history_disabled = 1;
                            selected_item = 0;
                            selected = 0;
                        end
                    end
                endcase
                // ǥ�õǴ� ���� �� �ݾ� ������ ���� �ֱ� ������ ����
                display_money_binary = total_money_history[7*9-1:7*8];
            end
            else if (return_sw) begin
                // ǥ�õǴ� ���� �� �ݾ� ������ ���� �ֱ� ������ ����
                display_money_binary = total_money_history[7*9-1:7*8];
                // return state Ȱ��ȭ
                return_state = 1;
            end

            // fnd array�� ���� if�� ��

            // ���� �Է� ��ư�� �������� ��
            if (coin_btn_state) begin
                // ǥ�õ� cnt���� �Ѿ��� ��
                if (coin_btn_cnt >= coin_btn_cnt_limit) begin
                    coin_btn_cnt = 0;
                    coin_btn_state = 0;
                    // ǥ�õǴ� ���� �� �ݾ� ������ ���� �ֱ� ������ �ǵ��� ��
                    display_money_binary = total_money_history[7*9-1:7*8];
                end 
                else coin_btn_cnt = coin_btn_cnt + 1;
            end
            // ��ȯ ��ư�� �������� ��
            else if (return_state) begin
                if (return_cnt >= return_cnt_limit) begin
                    return_cnt = 0;
                    // ���� ���°� �ƴ� ��
                    if (!history_disabled) begin
                        // �� �ݾ� ���縦 �� �ܰ辿 ������ �ǵ��� ��
                        total_money_history[7*9-1:7*1] = total_money_history[7*8-1:7*0];
                        total_money_history[7*1-1:7*0] = 8'd0;
                        display_money_binary = total_money_history[7*9-1:7*8];
                        if (total_money_history == 0) return_state = 0;                 
                    end
                    else begin
                        // ���� ������ ��� �� �ݾ� ���� ���� �ֱ� �ݾ��� 1�� ����
                        // 100���� ��ȯ�Ǵ� ��� ����
                        if (total_money_history[7*9-1:7*8] != 0) begin
                            total_money_history[7*9-1:7*8] = total_money_history[7*9-1:7*8] - 1;
                            display_money_binary = total_money_history[7*9-1:7*8];
                        end
                        else begin
                            // �� �ݾ��� 0���� ���� �� return state ��ȿȭ
                            return_state = 0;
                            history_disabled = 0;
                        end
                    end
                end
                else return_cnt = return_cnt + 1;
            end
            
            // lcd�� ���� if��
            case (cursor_pos)
                0 : begin
                    // prod 1, prod 2
                    line1_prod = prod1_id;
                    line2_prod = prod2_id;
                end
                1 : begin
                    if (ddram_address == 7'h4d) begin
                        // prod 1, prod 2
                        line1_prod = prod1_id;
                        line2_prod = prod2_id;
                    end
                    else if (ddram_address == 7'hd) begin
                        // prod 2, prod 3
                        line1_prod = prod2_id;
                        line2_prod = prod3_id;
                    end
                end
                2 : begin
                    // prod 2, prod 3
                    line1_prod = prod2_id;
                    line2_prod = prod3_id;
                end
                default : begin
                    // prod 1, prod 2
                    line1_prod = prod1_id;
                    line2_prod = prod2_id;
                end
            endcase

            case (line1_prod)
                1 : begin
                    line1_text[8*16-1:8*9] = product[8*7*3-1:8*7*2];
                    line1_text[8*8-1:8*6] = price_text[8*2*3-1:8*2*2];
                    if (prod1_count == 0) line1_text[8*2-1:8*1] = 8'h58; // "X"
                    else line1_text[8*2-1:8*1] = 8'h20; // "space"

                    if (line1_prod == selected_item) line1_text[8*3-1:8*2] = 8'h2a; // "*"
                    else line1_text[8*3-1:8*2] = 8'h20; // space
                end
                2 : begin
                    line1_text[8*16-1:8*9] = product[8*7*2-1:8*7*1];
                    line1_text[8*8-1:8*6] = price_text[8*2*2-1:8*2*1];
                    if (prod2_count == 0) line1_text[8*2-1:8*1] = 8'h58; // "X"
                    else line1_text[8*2-1:8*1] = 8'h20; // "space"

                    if (line1_prod == selected_item) line1_text[8*3-1:8*2] = 8'h2a; // "*"
                    else line1_text[8*3-1:8*2] = 8'h20; // space
                end
                3 : begin
                    line1_text[8*16-1:8*9] = product[8*7*1-1:8*7*0];
                    line1_text[8*8-1:8*6] = price_text[8*2*1-1:8*2*0];
                    if (prod3_count == 0) line1_text[8*2-1:8*1] = 8'h58; // "X"
                    else line1_text[8*2-1:8*1] = 8'h20; // "space"

                    if (line1_prod == selected_item) line1_text[8*3-1:8*2] = 8'h2a; // "*"
                    else line1_text[8*3-1:8*2] = 8'h20; // space
                end
                default : begin
                    line1_text[8*16-1:8*9] = product[8*7*3-1:8*7*2];
                    line1_text[8*3-1:8*2] = 8'h20; // "space"
                    line1_text[8*2-1:8*1] = 8'h20; // "space"
                end
            endcase

            case (line2_prod)
                1 : begin
                    line2_text[8*16-1:8*9] = product[8*7*3-1:8*7*2];
                    line2_text[8*8-1:8*6] = price_text[8*2*3-1:8*2*2];
                    if (prod1_count == 0) line2_text[8*2-1:8*1] = 8'h58; // "X"
                    else line2_text[8*2-1:8*1] = 8'h20; // "space"
                
                    if (line2_prod == selected_item) line2_text[8*3-1:8*2] = 8'h2a; // "*"
                    else line2_text[8*3-1:8*2] = 8'h20; // space
                end
                2 : begin
                    line2_text[8*16-1:8*9] = product[8*7*2-1:8*7*1];
                    line2_text[8*8-1:8*6] = price_text[8*2*2-1:8*2*1];
                    if (prod2_count == 0) line2_text[8*2-1:8*1] = 8'h58; // "X"
                    else line2_text[8*2-1:8*1] = 8'h20; // "space"

                    if (line2_prod == selected_item) line2_text[8*3-1:8*2] = 8'h2a; // "*"
                    else line2_text[8*3-1:8*2] = 8'h20; // space
                end
                3 : begin
                    line2_text[8*16-1:8*9] = product[8*7*1-1:8*7*0];
                    line2_text[8*8-1:8*6] = price_text[8*2*1-1:8*2*0];
                    if (prod3_count == 0) line2_text[8*2-1:8*1] = 8'h58; // "X"
                    else line2_text[8*2-1:8*1] = 8'h20; // "space"

                    if (line2_prod == selected_item) line2_text[8*3-1:8*2] = 8'h2a; // "*"
                    else line2_text[8*3-1:8*2] = 8'h20; // space
                end
                default : begin
                    line2_text[8*16-1:8*9] = product[8*7*2-1:8*7*1];
                    line2_text[8*3-1:8*2] = 8'h20; // "space"
                    line2_text[8*2-1:8*1] = 8'h20; // "space"
                end
            endcase
        end
    end
endmodule
